library verilog;
use verilog.vl_types.all;
entity addsub_vlg_vec_tst is
end addsub_vlg_vec_tst;
