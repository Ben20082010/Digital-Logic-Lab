library verilog;
use verilog.vl_types.all;
entity fourbitadd_vlg_vec_tst is
end fourbitadd_vlg_vec_tst;
