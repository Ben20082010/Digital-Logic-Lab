library verilog;
use verilog.vl_types.all;
entity extALU_vlg_vec_tst is
end extALU_vlg_vec_tst;
