library verilog;
use verilog.vl_types.all;
entity Nand2sim_vlg_vec_tst is
end Nand2sim_vlg_vec_tst;
