library verilog;
use verilog.vl_types.all;
entity alutest_vlg_vec_tst is
end alutest_vlg_vec_tst;
